library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
library lattice;
use lattice.all;
library machxo2;
use machxo2.all;

use packagekey00.all;

entity key00 is
	port(
		cdiv0:in std_logic_vector(4 downto 0);
		en0:std_logic;
		inkey0:in std_logic_vector(3 downto 0);
		clk0:inout std_logic;
		outr0:out std_logic_vector(3 downto 0);
		outcoder0:out std_logic_vector(6 downto 0)
	);
end key00;

architecture key0 of key00 is
signal outr00:std_logic_vector(3 downto 0);
begin
	k00: osc00 port map(
						cdiv=>cdiv0,
						oscOut0=>clk0
					);

	k01: contring00 port map(
							clkr=>clk0,
							enr=>en0,
							outr=>outr00
						);

	k02: coder00 port map(
							clkc=>clk0,
							incontc=>outr00,
							inkeyc=>inkey0,
							outcoder=>outcoder0
						);
	outr0<=outr00;

end key0;