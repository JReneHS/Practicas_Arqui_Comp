library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library lattice;
use lattice.all;
library machxo2;
use machxo2.all;

entity memrom00 is
	port(
		clkm:in std_logic
	);
end memrom00;

architecture memrom0 of memrom00 is
begin
end memrom0;